library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
entity clk_wiz_0_clk_wiz_0_clk_wiz is
	port (
			 clk_in1 : in STD_LOGIC;
			 clk_out1 : out STD_LOGIC;
			 clk_out2 : out STD_LOGIC;
			 clk_out3 : out STD_LOGIC;
			 clk_out4 : out STD_LOGIC;
			 reset : in STD_LOGIC;
			 locked : out STD_LOGIC
		 );
	attribute ORIG_REF_NAME : string;
	attribute ORIG_REF_NAME of clk_wiz_0_clk_wiz_0_clk_wiz : entity is "clk_wiz_0_clk_wiz";
end clk_wiz_0_clk_wiz_0_clk_wiz;

architecture STRUCTURE of clk_wiz_0_clk_wiz_0_clk_wiz is
	signal clk_in1_clk_wiz_0 : STD_LOGIC;
	signal clk_out1_clk_wiz_0 : STD_LOGIC;
	signal clk_out2_clk_wiz_0 : STD_LOGIC;
	signal clk_out3_clk_wiz_0 : STD_LOGIC;
	signal clk_out4_clk_wiz_0 : STD_LOGIC;
	signal clkfbout_buf_clk_wiz_0 : STD_LOGIC;
	signal clkfbout_clk_wiz_0 : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKFBOUTB_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKFBSTOPPED_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKINSTOPPED_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT0B_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT1B_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT2B_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT3B_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT4_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT5_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_CLKOUT6_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_DRDY_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_PSDONE_UNCONNECTED : STD_LOGIC;
	signal NLW_mmcm_adv_inst_DO_UNCONNECTED : STD_LOGIC_VECTOR ( 15 downto 0 );
	attribute BOX_TYPE : string;
	attribute BOX_TYPE of clkf_buf : label is "PRIMITIVE";
	attribute BOX_TYPE of clkin1_ibufg : label is "PRIMITIVE";
	attribute CAPACITANCE : string;
	attribute CAPACITANCE of clkin1_ibufg : label is "DONT_CARE";
	attribute IBUF_DELAY_VALUE : string;
	attribute IBUF_DELAY_VALUE of clkin1_ibufg : label is "0";
	attribute IFD_DELAY_VALUE : string;
	attribute IFD_DELAY_VALUE of clkin1_ibufg : label is "AUTO";
	attribute BOX_TYPE of clkout1_buf : label is "PRIMITIVE";
	attribute BOX_TYPE of clkout2_buf : label is "PRIMITIVE";
	attribute BOX_TYPE of clkout3_buf : label is "PRIMITIVE";
	attribute BOX_TYPE of clkout4_buf : label is "PRIMITIVE";
	attribute BOX_TYPE of mmcm_adv_inst : label is "PRIMITIVE";
begin
	clkf_buf: unisim.vcomponents.BUFG
	port map (
				 I => clkfbout_clk_wiz_0,
				 O => clkfbout_buf_clk_wiz_0
			 );
	clkin1_ibufg: unisim.vcomponents.IBUF
	generic map(
				   IOSTANDARD => "DEFAULT"
			   )
	port map (
				 I => clk_in1,
				 O => clk_in1_clk_wiz_0
			 );
	clkout1_buf: unisim.vcomponents.BUFG
	port map (
				 I => clk_out1_clk_wiz_0,
				 O => clk_out1
			 );
	clkout2_buf: unisim.vcomponents.BUFG
	port map (
				 I => clk_out2_clk_wiz_0,
				 O => clk_out2
			 );
	clkout3_buf: unisim.vcomponents.BUFG
	port map (
				 I => clk_out3_clk_wiz_0,
				 O => clk_out3
			 );
	clkout4_buf: unisim.vcomponents.BUFG
	port map (
				 I => clk_out4_clk_wiz_0,
				 O => clk_out4
			 );
	mmcm_adv_inst: unisim.vcomponents.MMCME2_ADV
	generic map(
				   BANDWIDTH => "OPTIMIZED",
				   CLKFBOUT_MULT_F => 6.000000,
				   CLKFBOUT_PHASE => 0.000000,
				   CLKFBOUT_USE_FINE_PS => false,
				   CLKIN1_PERIOD => 10.000000,
				   CLKIN2_PERIOD => 0.000000,
				   CLKOUT0_DIVIDE_F => 6.000000,
				   CLKOUT0_DUTY_CYCLE => 0.500000,
				   CLKOUT0_PHASE => 0.000000,
				   CLKOUT0_USE_FINE_PS => false,
				   CLKOUT1_DIVIDE => 3,
				   CLKOUT1_DUTY_CYCLE => 0.500000,
				   CLKOUT1_PHASE => 0.000000,
				   CLKOUT1_USE_FINE_PS => false,
				   CLKOUT2_DIVIDE => 50,
				   CLKOUT2_DUTY_CYCLE => 0.500000,
				   CLKOUT2_PHASE => 0.000000,
				   CLKOUT2_USE_FINE_PS => false,
				   CLKOUT3_DIVIDE => 12,
				   CLKOUT3_DUTY_CYCLE => 0.500000,
				   CLKOUT3_PHASE => 0.000000,
				   CLKOUT3_USE_FINE_PS => false,
				   CLKOUT4_CASCADE => false,
				   CLKOUT4_DIVIDE => 1,
				   CLKOUT4_DUTY_CYCLE => 0.500000,
				   CLKOUT4_PHASE => 0.000000,
				   CLKOUT4_USE_FINE_PS => false,
				   CLKOUT5_DIVIDE => 1,
				   CLKOUT5_DUTY_CYCLE => 0.500000,
				   CLKOUT5_PHASE => 0.000000,
				   CLKOUT5_USE_FINE_PS => false,
				   CLKOUT6_DIVIDE => 1,
				   CLKOUT6_DUTY_CYCLE => 0.500000,
				   CLKOUT6_PHASE => 0.000000,
				   CLKOUT6_USE_FINE_PS => false,
				   COMPENSATION => "ZHOLD",
				   DIVCLK_DIVIDE => 1,
				   IS_CLKINSEL_INVERTED => '0',
				   IS_PSEN_INVERTED => '0',
				   IS_PSINCDEC_INVERTED => '0',
				   IS_PWRDWN_INVERTED => '0',
				   IS_RST_INVERTED => '0',
				   REF_JITTER1 => 0.010000,
				   REF_JITTER2 => 0.010000,
				   SS_EN => "FALSE",
				   SS_MODE => "CENTER_HIGH",
				   SS_MOD_PERIOD => 10000,
				   STARTUP_WAIT => false
			   )
	port map (
				 CLKFBIN => clkfbout_buf_clk_wiz_0,
				 CLKFBOUT => clkfbout_clk_wiz_0,
				 CLKFBOUTB => NLW_mmcm_adv_inst_CLKFBOUTB_UNCONNECTED,
				 CLKFBSTOPPED => NLW_mmcm_adv_inst_CLKFBSTOPPED_UNCONNECTED,
				 CLKIN1 => clk_in1_clk_wiz_0,
				 CLKIN2 => '0',
				 CLKINSEL => '1',
				 CLKINSTOPPED => NLW_mmcm_adv_inst_CLKINSTOPPED_UNCONNECTED,
				 CLKOUT0 => clk_out1_clk_wiz_0,
				 CLKOUT0B => NLW_mmcm_adv_inst_CLKOUT0B_UNCONNECTED,
				 CLKOUT1 => clk_out2_clk_wiz_0,
				 CLKOUT1B => NLW_mmcm_adv_inst_CLKOUT1B_UNCONNECTED,
				 CLKOUT2 => clk_out3_clk_wiz_0,
				 CLKOUT2B => NLW_mmcm_adv_inst_CLKOUT2B_UNCONNECTED,
				 CLKOUT3 => clk_out4_clk_wiz_0,
				 CLKOUT3B => NLW_mmcm_adv_inst_CLKOUT3B_UNCONNECTED,
				 CLKOUT4 => NLW_mmcm_adv_inst_CLKOUT4_UNCONNECTED,
				 CLKOUT5 => NLW_mmcm_adv_inst_CLKOUT5_UNCONNECTED,
				 CLKOUT6 => NLW_mmcm_adv_inst_CLKOUT6_UNCONNECTED,
				 DADDR(6 downto 0) => B"0000000",
				 DCLK => '0',
				 DEN => '0',
				 DI(15 downto 0) => B"0000000000000000",
				 DO(15 downto 0) => NLW_mmcm_adv_inst_DO_UNCONNECTED(15 downto 0),
				 DRDY => NLW_mmcm_adv_inst_DRDY_UNCONNECTED,
				 DWE => '0',
				 LOCKED => locked,
				 PSCLK => '0',
				 PSDONE => NLW_mmcm_adv_inst_PSDONE_UNCONNECTED,
				 PSEN => '0',
				 PSINCDEC => '0',
				 PWRDWN => '0',
				 RST => reset
			 );
end STRUCTURE;

